vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|10 Mar 2014 11:53:48 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|10 Mar 2014 11:53:48 -0000
vti_filesize:IR|463
vti_backlinkinfo:VX|
