vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|24 Sep 2013 19:50:33 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|24 Sep 2013 19:50:33 -0000
vti_filesize:IR|24703
vti_backlinkinfo:VX|
