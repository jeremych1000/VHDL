vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|04 Mar 2014 13:39:05 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|04 Mar 2014 13:39:05 -0000
vti_filesize:IR|1113
vti_backlinkinfo:VX|
