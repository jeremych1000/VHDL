vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|10 Sep 2013 09:27:55 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|10 Sep 2013 09:27:55 -0000
vti_filesize:IR|2278
vti_backlinkinfo:VX|
