vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|10 Sep 2013 09:30:17 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|10 Sep 2013 09:30:17 -0000
vti_filesize:IR|11624
vti_backlinkinfo:VX|
