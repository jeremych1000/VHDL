vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|14 Feb 2013 19:27:30 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|14 Feb 2013 19:27:30 -0000
vti_filesize:IR|1751
vti_backlinkinfo:VX|
