vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|01 Mar 2014 19:06:05 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|01 Mar 2014 19:06:05 -0000
vti_filesize:IR|1673
vti_backlinkinfo:VX|
