vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|14 Feb 2015 22:54:22 -0000
vti_extenderversion:SR|12.0.0.0
vti_backlinkinfo:VX|
vti_syncwith_localhost\\w\:\\vhdl/w\:/vhdl:TR|09 Sep 2011 22:16:12 -0000
vti_modifiedby:SR|IC\\tomcl
vti_author:SR|IC\\tomcl
vti_nexttolasttimemodified:TW|14 Feb 2015 22:54:16 -0000
vti_timecreated:TR|14 Feb 2015 22:54:22 -0000
vti_cacheddtm:TX|14 Feb 2015 22:54:16 -0000
vti_filesize:IR|2133
