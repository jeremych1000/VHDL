vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|07 Sep 2013 15:16:12 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|07 Sep 2013 15:16:12 -0000
vti_filesize:IR|6886
vti_backlinkinfo:VX|
