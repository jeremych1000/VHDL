vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|25 Sep 2013 15:13:52 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|25 Sep 2013 15:13:52 -0000
vti_filesize:IR|786
vti_backlinkinfo:VX|
