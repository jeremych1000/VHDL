vti_encoding:SR|utf8-nl
vti_timelastmodified:TR|01 Feb 2015 17:23:34 -0000
vti_extenderversion:SR|12.0.0.0
vti_cacheddtm:TX|09 Sep 2011 22:16:52 -0000
vti_filesize:IR|3673
vti_backlinkinfo:VX|
vti_syncwith_localhost\\w\:\\vhdl/w\:/vhdl:TR|09 Sep 2011 22:16:52 -0000
vti_modifiedby:SR|IC\\tomcl
